BZh91AY&SY�D4J s߀Ryg���������`�|�[Q����$���L��=O�i�@h&� 4 q�&�CM��ѦL@��h�L Ɏ2dшi����4ɈMi�1�L�140CF�1#	�M0�&H	�OSBi3�G�<�CM �&��� ��C���ͤ����#M�ƍ#��p���q{(�YLTCkE=���f�#pI��=��볧��m�`����չM���N9cDZ��]0����`[Pnj+�� �0rjQ�B�=�C�t�C}��� =��lX��W�]9�Oz���3X�L�h�I�C����*��b� �
�,2X��)�<�L�"0S[�P�~H��.���S��+�`4a�=�R���B�,(�
��ٖ#>�����h��,�e�UC	"���Ҥ�NqVWQ<�ٮ6Qwę�FM_�ݴC�0���6��	�����//t���+�+6�%P�|�P���#��`K �JD�V����b�'T�Y�T���HjA��9��ZA�7�77$1l�8R�ߺ��E��+	��QƁ����=�K������Y�d����I$�I'�F�h���Ϝ=Z�T����+���T�Cu\�ثH7�R��B�aF8Q%�2/���xV趃94���C�/�����Q1f1`���$�O��@��JH�Y4M!���ֻ!�!	��Ȇ&s��Ã���$A��p�+���O�!�K ��3�6��q��u��ڐ�,5�@P�Ä�DU�����6yql�*�\����-�]�'QS�w�:[��	m~`� w���P�F� ���+0w�ڵ�$���hq�u��0U���=&���fƍ�d��%>�I'�������ıj�A�c���r� �`�~�����o�f�6�j�R�������/�����*ݻF��S��*~���#�o��f�E�6l5����h^��fj1� ��ͷ��tJI���`�Y�2n�+�&�8�Uȸ��ّ�(�n֚1	 FƏSć<����NQ�3˷q��tf>��t�\��~�Ȉ���,ܻ�u݋+�`�BqP��;̩�d�!	=a"IŒ=
�fC	e���uHF&օ�^��(#gE5I�����ON����4��y�vϝ�ld;�:�K��\�K#CJ���їY�0ؤ�!vct�L���0;��)��(�}G_Wf��_;�A
QV� ۂ:��@�=�̆�OA�
��pѱF4 ğ&F`��Tj0��1�M� V��u<v�5�.��&I2t�j��Z��9�%��%���{``�vx,	8$&M����Y�] �9A�=�%y�����W��Σ�v�`&�������ヽ��� ��:����T!����H`�ڏ :M�kd���G_���/<�/��P�6}�p��U�����<�RB@,�w� �^�1b���`x=��Nä{����7�6�c8�!�cC��  l��'�{)�>6��A���6���xC�B�]{j^��S�%[�FXֵ�!%��2�����3��݂�������z���ϛ����������u��V(P�ˋ����1˿�d��."q�|�V�~�$��@T:�<�Q
��+\�j5��y��7I��9��31�9�Rs����K��÷��7s���5�y�w ,V.�p�!�h�