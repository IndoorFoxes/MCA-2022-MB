BZh91AY&SY��7� �ߌRxg����������  `?      "Gꁠ� � 2i�@�4 h8ɓF!���`��i�q�&�CL	��14�@�&M�&�L�bi��!�L�1M00&�#��M A"A �ɩ�	��ш5M4Dm&�MF�	&�a�
��C	1V������BZN�>{}���M�O��L������~�zn�2B����/(i�h�����ĤĈJ�C>$/sF����p�=�F,X�;���v��o.,��y�뷎p��JEl�U��JC��������B��A���d�vs63;����U0�]	<�ju##ĩ�ԥ3]����ԩ��bޝ�)�,��ɩP��h�����A���H��ѐ/�4^�zt#?/-y�1��N��P[<!��-�耛�hV{�B�̹0��d��DƁ�9؍ôh����Y��s����{�^�a��jtk$`��P,p�2%[K
��	Z�R�h�ŇYB����7`�y�m�H cp�cm�@	�a��t%ّ��]�?p�X�6L���Ð\3��f��VD���*z`��2�F%%#/$�aJIM��Q3cJ���-.W���hЦ���8j#x@��@b��_��u�R�4_�a�d#Vx B&N;R�  �?�#�K����B�Bq����E�t�B��>���Ń1P�5�w0̻���6q�,
T���%3yC�%����q��br�M��0.6������(�Iz@���� H��\��y���̪�oR7�5����#�a���m�ڑ����>?B3$Ai�6�:�ZKBD�86\�.�aKjS@M�^`5Z(<m��"y�<���c �dɓ�9�аG�-�l�;MIXc�D���2�N]\�gۉ2H�D���q"�	������A
U�`�R]�0*���܉��jS� �*23(�#v �jDk
�=B�bE@�.��^U`3���3z�S��q�Q=V�CΒ�ڎ�T��FD���Shp���^HcLi��i��c1 ���8Ra`�M#�Q���À\^�mo*�J�!�.��%ʱ\_6򥁬��\�h-���&��))�����Z/Z-�lIC��"{9�1]����G���-c`�K������hL0�%���(y8��3�Li�)
@�X�e Ma�kYh	�"J�H���	r������1!4I�'kzb�D�����V��V����P�J��.�W��
P#��çxxZ�|ǭ<��K��! ���MI�c Ǵ�S���X}��l=�&f�Y�b�����HQ�Òd!���p[o�.b�H�:���cA���*yd��q���H�j3_�l[
$��LLG�.01��������iq�:���ib��/(Z"��Ě�ȑҨ@^⨓S{N�]�aҒ��"��q$���8T�)�,�u���C	��%=�0�h��B���j䴍[:.�ZL̼,	��2h�>��̖��`x��a2�)i�0�:����4�FQ�����b���4����R��3�o�Ӱe&1�/Ș1��u�������"�(Hm��