BZh91AY&SY��2 +߀Ryg����������`�|�P(��(E $�z��@�   dɡ��рFa `&�4��q�&�#F	���h�#@1�L��M`&i�L� �%h����2�M&�$�&�@�ddښRB&�	�&���S�(�țH @iْIQB�94?��i!�$�D��#Մ�#�.SidJ.I=������s�{���~�d|�.��)BH��1k��5��!qI�u��RS��]F�v@/"�Dzq��] ���S]�߶��21����h���Z���l��由�,��+�TۏYz�ϞL�ز�&��+&�[g����*��W����N�d�^�q��5Z.�6�b_g�����9���=�8m�O�$���ްľAz^��A��.�9���(i����j�2�ζ����wz�)_���H،͔}���;�ٟ�R0��bl2�Tc齚l&J�1*���ަ��Q�V�W�g]�h�s6�;�e�̩�[�6t���-5����-8�ڭ�Lr��FW]���m]�F�M.ή���x��)�z���*��e����UUR��e�Q���<�wux��T�
�0�#!q{/݋T��Og)��	�</m�j{j٭�ٛo���۬j�ٝ�yI�%t�ɽi4�l��R��W�ئ��b�n��}j.�,�yё4����r��c���:�j������a��}&8��ؐ���6E�b' �p�;�d��Ӹ�x�G��8<�32�5h�137\c����c����Ֆ�{7��a����c���5��I��M61����'�x���3؅Q���,��q�xuqy����wMG{䙑�'�����S��g�iw��w��1:H�mU��6|���xL��ӛC�hZJ����c�qH�L�q1	����Y����Y)�>�m���fa�S�L�����c�mSMjU�U���Wc��n�hay.�T��zWe�[8Lc+�"�e��9��ةe��a��M���|bt�1�rX2�iɔ��~�s;������s|$��S���7�~�UE<��6ocy�:{s1<��C9�>��lwF��%��d����<��T�Jz&S�?���*e/<x���������h;���X���6�]ܔ�g>����k.���X�<���f�ta�N�iȯ;�T��e�I��N��H�(�u-ey9R%�x��v�B����A8�R�mor,%4�]��jm>~��i!�9X}l�i�ŕ-UQIO�R�R].T��Y%M۹N����^d�[��;rC�����Z��bV5e
����͖KAĭ���F��if��M6��(�k/dk#7�w�餅x���N����3�qJ���R�����c���Gã���7��I��}=]R�sn��Z)��	ۯ�x�����D�8�|�V�~^"��׽w)����U'VIZ))'��R,.Q����h�^S�b\ܟ�ؒo9�P�o,%��YC�딩���g0ZF��r��17(q�����	F�Yy��>,�r��U_�k������vd(��3��`��rG�c����H�'5Gct��|�y�aѩ�Ĝy1�shF�9IC���Y=Q�];S�Bw���noNòK�3�M��9�]�&�)Q5�E�Ώ+Y�����;:�����0R��vN�F��rE8P���2